`timescale 1ns/1ps

//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:    
// Design Name:
// Module Name:    alu
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

module alu_top(
               src1,       //1 bit source 1 (input)
               src2,       //1 bit source 2 (input)
               less,       //1 bit less     (input)
               A_invert,   //1 bit A_invert (input)
               B_invert,   //1 bit B_invert (input)
               cin,        //1 bit carry in (input)
               operation,  //operation      (input)
               result,     //1 bit result   (output)
               cout       //1 bit carry out(output)
               );

input         src1;
input         src2;
input         less;
input         A_invert;
input         B_invert;
input         cin;
input [2-1:0] operation;

output        result;
output        cout;

reg           result;

wire A, B, AND, OR, ADD;

// invert gate for input
assign A = src1 ^ A_invert;
assign B = src2 ^ B_invert;
assign AND = A & B;
assign OR = A | B;

// self-define adder.v
adder e1(
    .a (A),
    .b (B),
    .c_in (cin),
    .sum (ADD),
    .c_out(cout)
);

// operations
always@(*)
begin
    case(operation)
        2'b00: result = AND;
        2'b01: result = OR;
        2'b10: result = ADD;
        2'b11: result = less;
    endcase
end

endmodule
